-- Elementos de Sistemas
-- by Luciano Soares
-- comparador16.vhd

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.all;

entity comparador16 is
   port(
	     a    : in STD_LOGIC_VECTOR(15 downto 0);
       zr   : out STD_LOGIC;
       ng   : out STD_LOGIC
   );
end comparador16;

architecture rtl of comparador16 is
  -- Aqui declaramos sinais (fios auxiliares)
  -- e componentes (outros módulos) que serao
  -- utilizados nesse modulo.

begin
  -- Implementação vem aqui!

  zr <= '1' when a = "0000000000000000" else '0';

  --ng <= '1' when to_integer(signed(a)) <  0 else '0';
  
  ng <= '1' when a(15) = '1' else '0';

end architecture;
